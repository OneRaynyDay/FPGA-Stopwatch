module nexys3(
	
);

clocks clocks_ (// Outputs
				// TODO
				// Inputs
				// TODO
				);

counter counter_ (// Outputs
				// TODO
				// Inputs
				// TODO
				);

display display_ (// Outputs
				// TODO
				// Inputs
				// TODO
				);

endmodule
